module SimpleCPU (
    //Ports definition
    input logic clk,
    input logic reset,
    
);
    
endmodule