module ALU (

    //Port definition
    input logic [7:0] A,
    input logic [7:0] B,
    input logic [2:0] Cntr,
    output logic [2:0] ALUFlags,s
    output logic [7:0] R
);

//Parameters


//Signals


endmodule